`define ENABLE_SUPER_RES 1
// `define ENABLE_WS2812 1
