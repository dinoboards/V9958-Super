`define ENABLE_SUPER_RES 1
