// File src/palette.vhd translated with vhd2vl 3.0 VHDL to Verilog RTL translator
// vhd2vl settings:
//  * Verilog Module Declaration Style: 2001

// vhd2vl is Free (libre) Software:
//   Copyright (C) 2001-2023 Vincenzo Liguori - Ocean Logic Pty Ltd
//     http://www.ocean-logic.com
//   Modifications Copyright (C) 2006 Mark Gonzales - PMC Sierra Inc
//   Modifications (C) 2010 Shankar Giri
//   Modifications Copyright (C) 2002-2023 Larry Doolittle
//     http://doolittle.icarus.com/~larry/vhd2vl/
//   Modifications (C) 2017 Rodrigo A. Melo
//
//   vhd2vl comes with ABSOLUTELY NO WARRANTY.  Always check the resulting
//   Verilog for correctness, ideally with a formal verification tool.
//
//   You are welcome to redistribute vhd2vl under certain conditions.
//   See the license (GPLv2) file included with the source for details.

// The result of translation follows.  Its copyright status should be
// considered unchanged from the original VHDL.

module PALETTE_RB (
    input wire [7:0] ADR,
    input wire CLK,
    input wire WE,
    input wire [7:0] DBO,
    output wire [7:0] DBI
);

  reg [7:0] blkram[0:255] = '{
      8'h00,
      8'h00,
      8'h11,
      8'h33,
      8'h26,
      8'h37,
      8'h52,
      8'h27,
      8'h62,
      8'h63,
      8'h52,
      8'h63,
      8'h11,
      8'h55,
      8'h55,
      8'h77,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00,
      8'h00
  };
  reg [7:0] iadr;

  always @(posedge CLK) begin
    if ((WE == 1'b1)) begin
      blkram[ADR] <= DBO;
    end
    iadr <= ADR;
  end

  assign DBI = blkram[iadr];

endmodule
