`define LEFT_BORDER 255

`define OFFSET_X 7'b0110101 // 49
`define LED_TV_X_NTSC  -20
`define LED_TV_Y_NTSC  1
`define LED_TV_X_PAL  -20
`define LED_TV_Y_PAL  3
